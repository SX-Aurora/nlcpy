global-exclude *.o *.c *.h *.cpp *.pyx *.pxi *.m4 *.master *.master2
include nlcpy/include/*.h
include nlcpy/veo/*.pxd
